// 64-bit ALU test bench template
module alu64bit_test;

// Put your code here
// ------------------


// End of your code

endmodule
